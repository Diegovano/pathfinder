// nio2_sys_tb.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module nio2_sys_tb (
	);

	wire         nio2_sys_inst_clk_bfm_clk_clk;       // nio2_sys_inst_clk_bfm:clk -> [nio2_sys_inst:clk_clk, nio2_sys_inst_reset_bfm:clk, sdram_my_partner:clk]
	wire         nio2_sys_inst_sdram_wire_cs_n;       // nio2_sys_inst:sdram_wire_cs_n -> sdram_my_partner:zs_cs_n
	wire   [1:0] nio2_sys_inst_sdram_wire_dqm;        // nio2_sys_inst:sdram_wire_dqm -> sdram_my_partner:zs_dqm
	wire         nio2_sys_inst_sdram_wire_cas_n;      // nio2_sys_inst:sdram_wire_cas_n -> sdram_my_partner:zs_cas_n
	wire         nio2_sys_inst_sdram_wire_ras_n;      // nio2_sys_inst:sdram_wire_ras_n -> sdram_my_partner:zs_ras_n
	wire         nio2_sys_inst_sdram_wire_we_n;       // nio2_sys_inst:sdram_wire_we_n -> sdram_my_partner:zs_we_n
	wire  [11:0] nio2_sys_inst_sdram_wire_addr;       // nio2_sys_inst:sdram_wire_addr -> sdram_my_partner:zs_addr
	wire         nio2_sys_inst_sdram_wire_cke;        // nio2_sys_inst:sdram_wire_cke -> sdram_my_partner:zs_cke
	wire  [15:0] nio2_sys_inst_sdram_wire_dq;         // [] -> [nio2_sys_inst:sdram_wire_dq, sdram_my_partner:zs_dq]
	wire   [1:0] nio2_sys_inst_sdram_wire_ba;         // nio2_sys_inst:sdram_wire_ba -> sdram_my_partner:zs_ba
	wire         nio2_sys_inst_reset_bfm_reset_reset; // nio2_sys_inst_reset_bfm:reset -> nio2_sys_inst:reset_reset_n

	nio2_sys nio2_sys_inst (
		.clk_clk                            (nio2_sys_inst_clk_bfm_clk_clk),       //                         clk.clk
		.led_pio_external_connection_export (),                                    // led_pio_external_connection.export
		.reset_reset_n                      (nio2_sys_inst_reset_bfm_reset_reset), //                       reset.reset_n
		.sdram_wire_addr                    (nio2_sys_inst_sdram_wire_addr),       //                  sdram_wire.addr
		.sdram_wire_ba                      (nio2_sys_inst_sdram_wire_ba),         //                            .ba
		.sdram_wire_cas_n                   (nio2_sys_inst_sdram_wire_cas_n),      //                            .cas_n
		.sdram_wire_cke                     (nio2_sys_inst_sdram_wire_cke),        //                            .cke
		.sdram_wire_cs_n                    (nio2_sys_inst_sdram_wire_cs_n),       //                            .cs_n
		.sdram_wire_dq                      (nio2_sys_inst_sdram_wire_dq),         //                            .dq
		.sdram_wire_dqm                     (nio2_sys_inst_sdram_wire_dqm),        //                            .dqm
		.sdram_wire_ras_n                   (nio2_sys_inst_sdram_wire_ras_n),      //                            .ras_n
		.sdram_wire_we_n                    (nio2_sys_inst_sdram_wire_we_n)        //                            .we_n
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) nio2_sys_inst_clk_bfm (
		.clk (nio2_sys_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) nio2_sys_inst_reset_bfm (
		.reset (nio2_sys_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (nio2_sys_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_sdram_partner_module sdram_my_partner (
		.clk      (nio2_sys_inst_clk_bfm_clk_clk),  //     clk.clk
		.zs_dq    (nio2_sys_inst_sdram_wire_dq),    // conduit.dq
		.zs_addr  (nio2_sys_inst_sdram_wire_addr),  //        .addr
		.zs_ba    (nio2_sys_inst_sdram_wire_ba),    //        .ba
		.zs_cas_n (nio2_sys_inst_sdram_wire_cas_n), //        .cas_n
		.zs_cke   (nio2_sys_inst_sdram_wire_cke),   //        .cke
		.zs_cs_n  (nio2_sys_inst_sdram_wire_cs_n),  //        .cs_n
		.zs_dqm   (nio2_sys_inst_sdram_wire_dqm),   //        .dqm
		.zs_ras_n (nio2_sys_inst_sdram_wire_ras_n), //        .ras_n
		.zs_we_n  (nio2_sys_inst_sdram_wire_we_n)   //        .we_n
	);

endmodule
